module top(
  input [7:0] a,
  input [7:0] b,
  input clk,
  input rst,
  output [15:0] led
  );
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_CE;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_I;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A0;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A1;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A10;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A11;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A12;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A13;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A14;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A15;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A16;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A17;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A18;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A19;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A2;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A20;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A21;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A22;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A23;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A24;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A25;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A26;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A27;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A28;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A29;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A3;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A4;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A5;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A6;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A7;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A8;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_A9;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT0;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT1;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT10;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT11;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT12;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT13;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT14;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT15;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT16;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT17;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT18;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT19;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT2;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT20;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT21;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT22;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT23;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT24;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT25;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT26;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT27;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT28;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT29;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT3;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT4;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT5;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT6;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT7;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT8;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ACOUT9;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ALUMODE0;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ALUMODE1;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ALUMODE2;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_ALUMODE3;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_B0;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_B1;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_B10;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_B11;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_B12;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_B13;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_B14;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_B15;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_B16;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_B17;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_B2;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_B3;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_B4;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_B5;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_B6;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_B7;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_B8;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_B9;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_BCOUT0;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_BCOUT1;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_BCOUT10;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_BCOUT11;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_BCOUT12;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_BCOUT13;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_BCOUT14;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_BCOUT15;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_BCOUT16;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_BCOUT17;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_BCOUT2;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_BCOUT3;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_BCOUT4;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_BCOUT5;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_BCOUT6;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_BCOUT7;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_BCOUT8;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_BCOUT9;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C0;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C1;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C10;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C11;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C12;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C13;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C14;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C15;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C16;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C17;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C18;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C19;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C2;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C20;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C21;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C22;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C23;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C24;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C25;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C26;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C27;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C28;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C29;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C3;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C30;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C31;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C32;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C33;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C34;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C35;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C36;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C37;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C38;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C39;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C4;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C40;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C41;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C42;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C43;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C44;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C45;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C46;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C47;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C5;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C6;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C7;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C8;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_C9;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_CARRYINSEL0;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_CARRYINSEL1;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_CARRYINSEL2;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_CARRYOUT0;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_CARRYOUT1;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_CARRYOUT2;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_CARRYOUT3;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_CEA1;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_CEA2;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_CEAD;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_CEALUMODE;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_CEB1;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_CEB2;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_CEC;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_CECARRYIN;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_CECTRL;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_CED;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_CEINMODE;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_CEM;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_CEP;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_CLK;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D0;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D1;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D10;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D11;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D12;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D13;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D14;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D15;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D16;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D17;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D18;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D19;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D2;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D20;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D21;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D22;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D23;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D24;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D3;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D4;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D5;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D6;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D7;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D8;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_D9;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_INMODE0;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_INMODE1;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_INMODE2;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_INMODE3;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_INMODE4;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_OPMODE0;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_OPMODE1;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_OPMODE2;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_OPMODE3;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_OPMODE4;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_OPMODE5;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_OPMODE6;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P0;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P1;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P10;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P11;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P12;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P13;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P14;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P15;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P16;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P17;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P18;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P19;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P2;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P20;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P21;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P22;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P23;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P24;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P25;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P26;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P27;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P28;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P29;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P3;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P30;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P31;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P32;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P33;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P34;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P35;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P36;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P37;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P38;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P39;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P4;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P40;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P41;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P42;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P43;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P44;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P45;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P46;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P47;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P5;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P6;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P7;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P8;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_P9;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT0;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT1;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT10;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT11;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT12;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT13;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT14;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT15;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT16;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT17;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT18;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT19;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT2;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT20;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT21;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT22;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT23;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT24;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT25;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT26;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT27;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT28;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT29;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT3;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT30;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT31;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT32;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT33;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT34;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT35;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT36;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT37;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT38;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT39;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT4;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT40;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT41;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT42;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT43;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT44;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT45;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT46;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT47;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT5;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT6;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT7;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT8;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_PCOUT9;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_RSTA;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_RSTALUMODE;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_RSTB;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_RSTC;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_RSTCTRL;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_RSTD;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_RSTINMODE;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_RSTM;
  wire [0:0] DSP_R_X9Y20_DSP48_X0Y8_RSTP;
  wire [0:0] LIOB33_SING_X0Y0_IOB_X0Y0_O;
  wire [0:0] LIOB33_X0Y11_IOB_X0Y11_I;
  wire [0:0] LIOB33_X0Y11_IOB_X0Y12_I;
  wire [0:0] LIOB33_X0Y13_IOB_X0Y13_I;
  wire [0:0] LIOB33_X0Y17_IOB_X0Y18_O;
  wire [0:0] LIOB33_X0Y19_IOB_X0Y19_O;
  wire [0:0] LIOB33_X0Y19_IOB_X0Y20_O;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y1_O;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y2_O;
  wire [0:0] LIOB33_X0Y3_IOB_X0Y3_O;
  wire [0:0] LIOB33_X0Y3_IOB_X0Y4_O;
  wire [0:0] LIOB33_X0Y43_IOB_X0Y43_O;
  wire [0:0] LIOB33_X0Y5_IOB_X0Y5_I;
  wire [0:0] LIOB33_X0Y5_IOB_X0Y6_I;
  wire [0:0] LIOB33_X0Y7_IOB_X0Y7_I;
  wire [0:0] LIOB33_X0Y7_IOB_X0Y8_I;
  wire [0:0] LIOB33_X0Y9_IOB_X0Y10_I;
  wire [0:0] LIOB33_X0Y9_IOB_X0Y9_I;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_D1;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_OQ;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_T1;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_O;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_D;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_O;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y12_D;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y12_O;
  wire [0:0] LIOI3_X0Y17_OLOGIC_X0Y18_D1;
  wire [0:0] LIOI3_X0Y17_OLOGIC_X0Y18_OQ;
  wire [0:0] LIOI3_X0Y17_OLOGIC_X0Y18_T1;
  wire [0:0] LIOI3_X0Y17_OLOGIC_X0Y18_TQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_D1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_OQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_T1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_TQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_D1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_OQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_T1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_TQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_D1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_OQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_T1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_TQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_D1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_OQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_T1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_TQ;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y5_D;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y5_O;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y6_D;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y6_O;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y10_D;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y10_O;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y9_D;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y9_O;
  wire [0:0] RIOB33_X43Y25_IOB_X1Y26_I;
  wire [0:0] RIOB33_X43Y31_IOB_X1Y32_O;
  wire [0:0] RIOB33_X43Y37_IOB_X1Y37_O;
  wire [0:0] RIOB33_X43Y37_IOB_X1Y38_O;
  wire [0:0] RIOB33_X43Y39_IOB_X1Y39_I;
  wire [0:0] RIOB33_X43Y39_IOB_X1Y40_I;
  wire [0:0] RIOB33_X43Y43_IOB_X1Y43_I;
  wire [0:0] RIOB33_X43Y43_IOB_X1Y44_I;
  wire [0:0] RIOB33_X43Y45_IOB_X1Y45_I;
  wire [0:0] RIOB33_X43Y45_IOB_X1Y46_I;
  wire [0:0] RIOB33_X43Y47_IOB_X1Y47_I;
  wire [0:0] RIOB33_X43Y47_IOB_X1Y48_I;
  wire [0:0] RIOB33_X43Y61_IOB_X1Y61_O;
  wire [0:0] RIOB33_X43Y75_IOB_X1Y75_O;
  wire [0:0] RIOB33_X43Y75_IOB_X1Y76_O;
  wire [0:0] RIOB33_X43Y87_IOB_X1Y87_O;
  wire [0:0] RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_D1;
  wire [0:0] RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_OQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_T1;
  wire [0:0] RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_TQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y43_D;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y43_O;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y44_D;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y44_O;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_D1;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_OQ;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_T1;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_TQ;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_D1;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_OQ;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_T1;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_TQ;
  wire [0:0] RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_D1;
  wire [0:0] RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_OQ;
  wire [0:0] RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_T1;
  wire [0:0] RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_TQ;
  wire [0:0] RIOI3_X43Y25_ILOGIC_X1Y26_D;
  wire [0:0] RIOI3_X43Y25_ILOGIC_X1Y26_O;
  wire [0:0] RIOI3_X43Y39_ILOGIC_X1Y39_D;
  wire [0:0] RIOI3_X43Y39_ILOGIC_X1Y39_O;
  wire [0:0] RIOI3_X43Y39_ILOGIC_X1Y40_D;
  wire [0:0] RIOI3_X43Y39_ILOGIC_X1Y40_O;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y45_D;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y45_O;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y46_D;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y46_O;
  wire [0:0] RIOI3_X43Y47_ILOGIC_X1Y47_D;
  wire [0:0] RIOI3_X43Y47_ILOGIC_X1Y47_O;
  wire [0:0] RIOI3_X43Y47_ILOGIC_X1Y48_D;
  wire [0:0] RIOI3_X43Y47_ILOGIC_X1Y48_O;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_D1;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_OQ;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_T1;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_TQ;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y75_D1;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y75_OQ;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y75_T1;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y75_TQ;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y76_D1;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y76_OQ;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y76_T1;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y76_TQ;


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(RIOB33_X43Y25_IOB_X1Y26_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "DSP48E1" *)
  DSP48E1 #(
    .ACASCREG(1),
    .AREG(1),
    .A_INPUT("DIRECT"),
    .BCASCREG(1),
    .BREG(1),
    .B_INPUT("DIRECT")
  ) DSP_R_X9Y20_DSP48_X0Y8_DSP48E1 (
.A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, LIOB33_X0Y5_IOB_X0Y6_I, LIOB33_X0Y5_IOB_X0Y5_I, LIOB33_X0Y7_IOB_X0Y8_I, LIOB33_X0Y7_IOB_X0Y7_I, LIOB33_X0Y9_IOB_X0Y9_I, LIOB33_X0Y9_IOB_X0Y10_I, LIOB33_X0Y11_IOB_X0Y12_I, LIOB33_X0Y11_IOB_X0Y11_I}),
.ACOUT({DSP_R_X9Y20_DSP48_X0Y8_ACOUT29, DSP_R_X9Y20_DSP48_X0Y8_ACOUT28, DSP_R_X9Y20_DSP48_X0Y8_ACOUT27, DSP_R_X9Y20_DSP48_X0Y8_ACOUT26, DSP_R_X9Y20_DSP48_X0Y8_ACOUT25, DSP_R_X9Y20_DSP48_X0Y8_ACOUT24, DSP_R_X9Y20_DSP48_X0Y8_ACOUT23, DSP_R_X9Y20_DSP48_X0Y8_ACOUT22, DSP_R_X9Y20_DSP48_X0Y8_ACOUT21, DSP_R_X9Y20_DSP48_X0Y8_ACOUT20, DSP_R_X9Y20_DSP48_X0Y8_ACOUT19, DSP_R_X9Y20_DSP48_X0Y8_ACOUT18, DSP_R_X9Y20_DSP48_X0Y8_ACOUT17, DSP_R_X9Y20_DSP48_X0Y8_ACOUT16, DSP_R_X9Y20_DSP48_X0Y8_ACOUT15, DSP_R_X9Y20_DSP48_X0Y8_ACOUT14, DSP_R_X9Y20_DSP48_X0Y8_ACOUT13, DSP_R_X9Y20_DSP48_X0Y8_ACOUT12, DSP_R_X9Y20_DSP48_X0Y8_ACOUT11, DSP_R_X9Y20_DSP48_X0Y8_ACOUT10, DSP_R_X9Y20_DSP48_X0Y8_ACOUT9, DSP_R_X9Y20_DSP48_X0Y8_ACOUT8, DSP_R_X9Y20_DSP48_X0Y8_ACOUT7, DSP_R_X9Y20_DSP48_X0Y8_ACOUT6, DSP_R_X9Y20_DSP48_X0Y8_ACOUT5, DSP_R_X9Y20_DSP48_X0Y8_ACOUT4, DSP_R_X9Y20_DSP48_X0Y8_ACOUT3, DSP_R_X9Y20_DSP48_X0Y8_ACOUT2, DSP_R_X9Y20_DSP48_X0Y8_ACOUT1, DSP_R_X9Y20_DSP48_X0Y8_ACOUT0}),
.ALUMODE({1'b0, 1'b0, 1'b1, 1'b1}),
.B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, RIOB33_X43Y47_IOB_X1Y48_I, RIOB33_X43Y43_IOB_X1Y44_I, RIOB33_X43Y43_IOB_X1Y43_I, RIOB33_X43Y39_IOB_X1Y39_I, RIOB33_X43Y45_IOB_X1Y46_I, RIOB33_X43Y47_IOB_X1Y47_I, RIOB33_X43Y45_IOB_X1Y45_I, RIOB33_X43Y39_IOB_X1Y40_I}),
.BCOUT({DSP_R_X9Y20_DSP48_X0Y8_BCOUT17, DSP_R_X9Y20_DSP48_X0Y8_BCOUT16, DSP_R_X9Y20_DSP48_X0Y8_BCOUT15, DSP_R_X9Y20_DSP48_X0Y8_BCOUT14, DSP_R_X9Y20_DSP48_X0Y8_BCOUT13, DSP_R_X9Y20_DSP48_X0Y8_BCOUT12, DSP_R_X9Y20_DSP48_X0Y8_BCOUT11, DSP_R_X9Y20_DSP48_X0Y8_BCOUT10, DSP_R_X9Y20_DSP48_X0Y8_BCOUT9, DSP_R_X9Y20_DSP48_X0Y8_BCOUT8, DSP_R_X9Y20_DSP48_X0Y8_BCOUT7, DSP_R_X9Y20_DSP48_X0Y8_BCOUT6, DSP_R_X9Y20_DSP48_X0Y8_BCOUT5, DSP_R_X9Y20_DSP48_X0Y8_BCOUT4, DSP_R_X9Y20_DSP48_X0Y8_BCOUT3, DSP_R_X9Y20_DSP48_X0Y8_BCOUT2, DSP_R_X9Y20_DSP48_X0Y8_BCOUT1, DSP_R_X9Y20_DSP48_X0Y8_BCOUT0}),
.C({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.CARRYINSEL({1'b0, 1'b0, 1'b0}),
.CARRYOUT({DSP_R_X9Y20_DSP48_X0Y8_CARRYOUT3, DSP_R_X9Y20_DSP48_X0Y8_CARRYOUT2, DSP_R_X9Y20_DSP48_X0Y8_CARRYOUT1, DSP_R_X9Y20_DSP48_X0Y8_CARRYOUT0}),
.CEA1(1'b0),
.CEA2(1'b1),
.CEAD(1'b0),
.CEALUMODE(1'b0),
.CEB1(1'b0),
.CEB2(1'b1),
.CEC(1'b0),
.CECARRYIN(1'b0),
.CECTRL(1'b0),
.CED(1'b0),
.CEINMODE(1'b0),
.CEM(1'b1),
.CEP(1'b1),
.CLK(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.D({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.INMODE({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.OPMODE({1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.P({DSP_R_X9Y20_DSP48_X0Y8_P47, DSP_R_X9Y20_DSP48_X0Y8_P46, DSP_R_X9Y20_DSP48_X0Y8_P45, DSP_R_X9Y20_DSP48_X0Y8_P44, DSP_R_X9Y20_DSP48_X0Y8_P43, DSP_R_X9Y20_DSP48_X0Y8_P42, DSP_R_X9Y20_DSP48_X0Y8_P41, DSP_R_X9Y20_DSP48_X0Y8_P40, DSP_R_X9Y20_DSP48_X0Y8_P39, DSP_R_X9Y20_DSP48_X0Y8_P38, DSP_R_X9Y20_DSP48_X0Y8_P37, DSP_R_X9Y20_DSP48_X0Y8_P36, DSP_R_X9Y20_DSP48_X0Y8_P35, DSP_R_X9Y20_DSP48_X0Y8_P34, DSP_R_X9Y20_DSP48_X0Y8_P33, DSP_R_X9Y20_DSP48_X0Y8_P32, DSP_R_X9Y20_DSP48_X0Y8_P31, DSP_R_X9Y20_DSP48_X0Y8_P30, DSP_R_X9Y20_DSP48_X0Y8_P29, DSP_R_X9Y20_DSP48_X0Y8_P28, DSP_R_X9Y20_DSP48_X0Y8_P27, DSP_R_X9Y20_DSP48_X0Y8_P26, DSP_R_X9Y20_DSP48_X0Y8_P25, DSP_R_X9Y20_DSP48_X0Y8_P24, DSP_R_X9Y20_DSP48_X0Y8_P23, DSP_R_X9Y20_DSP48_X0Y8_P22, DSP_R_X9Y20_DSP48_X0Y8_P21, DSP_R_X9Y20_DSP48_X0Y8_P20, DSP_R_X9Y20_DSP48_X0Y8_P19, DSP_R_X9Y20_DSP48_X0Y8_P18, DSP_R_X9Y20_DSP48_X0Y8_P17, DSP_R_X9Y20_DSP48_X0Y8_P16, DSP_R_X9Y20_DSP48_X0Y8_P15, DSP_R_X9Y20_DSP48_X0Y8_P14, DSP_R_X9Y20_DSP48_X0Y8_P13, DSP_R_X9Y20_DSP48_X0Y8_P12, DSP_R_X9Y20_DSP48_X0Y8_P11, DSP_R_X9Y20_DSP48_X0Y8_P10, DSP_R_X9Y20_DSP48_X0Y8_P9, DSP_R_X9Y20_DSP48_X0Y8_P8, DSP_R_X9Y20_DSP48_X0Y8_P7, DSP_R_X9Y20_DSP48_X0Y8_P6, DSP_R_X9Y20_DSP48_X0Y8_P5, DSP_R_X9Y20_DSP48_X0Y8_P4, DSP_R_X9Y20_DSP48_X0Y8_P3, DSP_R_X9Y20_DSP48_X0Y8_P2, DSP_R_X9Y20_DSP48_X0Y8_P1, DSP_R_X9Y20_DSP48_X0Y8_P0}),
.PCOUT({DSP_R_X9Y20_DSP48_X0Y8_PCOUT47, DSP_R_X9Y20_DSP48_X0Y8_PCOUT46, DSP_R_X9Y20_DSP48_X0Y8_PCOUT45, DSP_R_X9Y20_DSP48_X0Y8_PCOUT44, DSP_R_X9Y20_DSP48_X0Y8_PCOUT43, DSP_R_X9Y20_DSP48_X0Y8_PCOUT42, DSP_R_X9Y20_DSP48_X0Y8_PCOUT41, DSP_R_X9Y20_DSP48_X0Y8_PCOUT40, DSP_R_X9Y20_DSP48_X0Y8_PCOUT39, DSP_R_X9Y20_DSP48_X0Y8_PCOUT38, DSP_R_X9Y20_DSP48_X0Y8_PCOUT37, DSP_R_X9Y20_DSP48_X0Y8_PCOUT36, DSP_R_X9Y20_DSP48_X0Y8_PCOUT35, DSP_R_X9Y20_DSP48_X0Y8_PCOUT34, DSP_R_X9Y20_DSP48_X0Y8_PCOUT33, DSP_R_X9Y20_DSP48_X0Y8_PCOUT32, DSP_R_X9Y20_DSP48_X0Y8_PCOUT31, DSP_R_X9Y20_DSP48_X0Y8_PCOUT30, DSP_R_X9Y20_DSP48_X0Y8_PCOUT29, DSP_R_X9Y20_DSP48_X0Y8_PCOUT28, DSP_R_X9Y20_DSP48_X0Y8_PCOUT27, DSP_R_X9Y20_DSP48_X0Y8_PCOUT26, DSP_R_X9Y20_DSP48_X0Y8_PCOUT25, DSP_R_X9Y20_DSP48_X0Y8_PCOUT24, DSP_R_X9Y20_DSP48_X0Y8_PCOUT23, DSP_R_X9Y20_DSP48_X0Y8_PCOUT22, DSP_R_X9Y20_DSP48_X0Y8_PCOUT21, DSP_R_X9Y20_DSP48_X0Y8_PCOUT20, DSP_R_X9Y20_DSP48_X0Y8_PCOUT19, DSP_R_X9Y20_DSP48_X0Y8_PCOUT18, DSP_R_X9Y20_DSP48_X0Y8_PCOUT17, DSP_R_X9Y20_DSP48_X0Y8_PCOUT16, DSP_R_X9Y20_DSP48_X0Y8_PCOUT15, DSP_R_X9Y20_DSP48_X0Y8_PCOUT14, DSP_R_X9Y20_DSP48_X0Y8_PCOUT13, DSP_R_X9Y20_DSP48_X0Y8_PCOUT12, DSP_R_X9Y20_DSP48_X0Y8_PCOUT11, DSP_R_X9Y20_DSP48_X0Y8_PCOUT10, DSP_R_X9Y20_DSP48_X0Y8_PCOUT9, DSP_R_X9Y20_DSP48_X0Y8_PCOUT8, DSP_R_X9Y20_DSP48_X0Y8_PCOUT7, DSP_R_X9Y20_DSP48_X0Y8_PCOUT6, DSP_R_X9Y20_DSP48_X0Y8_PCOUT5, DSP_R_X9Y20_DSP48_X0Y8_PCOUT4, DSP_R_X9Y20_DSP48_X0Y8_PCOUT3, DSP_R_X9Y20_DSP48_X0Y8_PCOUT2, DSP_R_X9Y20_DSP48_X0Y8_PCOUT1, DSP_R_X9Y20_DSP48_X0Y8_PCOUT0}),
.RSTA(LIOB33_X0Y13_IOB_X0Y13_I),
.RSTALUMODE(1'b0),
.RSTB(LIOB33_X0Y13_IOB_X0Y13_I),
.RSTC(1'b0),
.RSTCTRL(1'b0),
.RSTD(1'b0),
.RSTINMODE(1'b0),
.RSTM(LIOB33_X0Y13_IOB_X0Y13_I),
.RSTP(LIOB33_X0Y13_IOB_X0Y13_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y1_IOB_X0Y1_OBUF (
.I(DSP_R_X9Y20_DSP48_X0Y8_P7),
.O(led[7])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y1_IOB_X0Y2_OBUF (
.I(DSP_R_X9Y20_DSP48_X0Y8_P8),
.O(led[8])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y3_IOB_X0Y3_OBUF (
.I(DSP_R_X9Y20_DSP48_X0Y8_P0),
.O(led[0])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y3_IOB_X0Y4_OBUF (
.I(DSP_R_X9Y20_DSP48_X0Y8_P5),
.O(led[5])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y5_IOB_X0Y5_IBUF (
.I(a[6]),
.O(LIOB33_X0Y5_IOB_X0Y5_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y5_IOB_X0Y6_IBUF (
.I(a[7]),
.O(LIOB33_X0Y5_IOB_X0Y6_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y7_IOB_X0Y7_IBUF (
.I(a[4]),
.O(LIOB33_X0Y7_IOB_X0Y7_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y7_IOB_X0Y8_IBUF (
.I(a[5]),
.O(LIOB33_X0Y7_IOB_X0Y8_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y9_IOB_X0Y9_IBUF (
.I(a[3]),
.O(LIOB33_X0Y9_IOB_X0Y9_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y9_IOB_X0Y10_IBUF (
.I(a[2]),
.O(LIOB33_X0Y9_IOB_X0Y10_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y11_IOB_X0Y11_IBUF (
.I(a[0]),
.O(LIOB33_X0Y11_IOB_X0Y11_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y11_IOB_X0Y12_IBUF (
.I(a[1]),
.O(LIOB33_X0Y11_IOB_X0Y12_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y13_IOB_X0Y13_IBUF (
.I(rst),
.O(LIOB33_X0Y13_IOB_X0Y13_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y17_IOB_X0Y18_OBUF (
.I(DSP_R_X9Y20_DSP48_X0Y8_P4),
.O(led[4])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y19_IOB_X0Y19_OBUF (
.I(DSP_R_X9Y20_DSP48_X0Y8_P3),
.O(led[3])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y19_IOB_X0Y20_OBUF (
.I(DSP_R_X9Y20_DSP48_X0Y8_P2),
.O(led[2])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y43_IOB_X0Y43_OBUF (
.I(DSP_R_X9Y20_DSP48_X0Y8_P1),
.O(led[1])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y0_IOB_X0Y0_OBUF (
.I(DSP_R_X9Y20_DSP48_X0Y8_P6),
.O(led[6])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X43Y25_IOB_X1Y26_IBUF (
.I(clk),
.O(RIOB33_X43Y25_IOB_X1Y26_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X43Y31_IOB_X1Y32_OBUF (
.I(DSP_R_X9Y20_DSP48_X0Y8_P11),
.O(led[11])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X43Y37_IOB_X1Y37_OBUF (
.I(DSP_R_X9Y20_DSP48_X0Y8_P10),
.O(led[10])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X43Y37_IOB_X1Y38_OBUF (
.I(DSP_R_X9Y20_DSP48_X0Y8_P9),
.O(led[9])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X43Y39_IOB_X1Y39_IBUF (
.I(b[4]),
.O(RIOB33_X43Y39_IOB_X1Y39_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X43Y39_IOB_X1Y40_IBUF (
.I(b[0]),
.O(RIOB33_X43Y39_IOB_X1Y40_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X43Y43_IOB_X1Y43_IBUF (
.I(b[5]),
.O(RIOB33_X43Y43_IOB_X1Y43_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X43Y43_IOB_X1Y44_IBUF (
.I(b[6]),
.O(RIOB33_X43Y43_IOB_X1Y44_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X43Y45_IOB_X1Y45_IBUF (
.I(b[1]),
.O(RIOB33_X43Y45_IOB_X1Y45_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X43Y45_IOB_X1Y46_IBUF (
.I(b[3]),
.O(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X43Y47_IOB_X1Y47_IBUF (
.I(b[2]),
.O(RIOB33_X43Y47_IOB_X1Y47_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X43Y47_IOB_X1Y48_IBUF (
.I(b[7]),
.O(RIOB33_X43Y47_IOB_X1Y48_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X43Y61_IOB_X1Y61_OBUF (
.I(DSP_R_X9Y20_DSP48_X0Y8_P14),
.O(led[14])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X43Y75_IOB_X1Y75_OBUF (
.I(DSP_R_X9Y20_DSP48_X0Y8_P12),
.O(led[12])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X43Y75_IOB_X1Y76_OBUF (
.I(DSP_R_X9Y20_DSP48_X0Y8_P13),
.O(led[13])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X43Y87_IOB_X1Y87_OBUF (
.I(DSP_R_X9Y20_DSP48_X0Y8_P15),
.O(led[15])
  );
  assign LIOI3_X0Y1_OLOGIC_X0Y2_OQ = DSP_R_X9Y20_DSP48_X0Y8_P8;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_TQ = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_OQ = DSP_R_X9Y20_DSP48_X0Y8_P7;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_TQ = 1'b1;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_OQ = DSP_R_X9Y20_DSP48_X0Y8_P5;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_TQ = 1'b1;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_OQ = DSP_R_X9Y20_DSP48_X0Y8_P0;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_TQ = 1'b1;
  assign LIOI3_X0Y5_ILOGIC_X0Y6_O = LIOB33_X0Y5_IOB_X0Y6_I;
  assign LIOI3_X0Y5_ILOGIC_X0Y5_O = LIOB33_X0Y5_IOB_X0Y5_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y10_O = LIOB33_X0Y9_IOB_X0Y10_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y9_O = LIOB33_X0Y9_IOB_X0Y9_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y12_O = LIOB33_X0Y11_IOB_X0Y12_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_O = LIOB33_X0Y11_IOB_X0Y11_I;
  assign LIOI3_X0Y17_OLOGIC_X0Y18_OQ = DSP_R_X9Y20_DSP48_X0Y8_P4;
  assign LIOI3_X0Y17_OLOGIC_X0Y18_TQ = 1'b1;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_OQ = DSP_R_X9Y20_DSP48_X0Y8_P6;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_O = LIOB33_X0Y7_IOB_X0Y8_I;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_O = LIOB33_X0Y7_IOB_X0Y7_I;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_OQ = DSP_R_X9Y20_DSP48_X0Y8_P2;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_OQ = DSP_R_X9Y20_DSP48_X0Y8_P3;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_OQ = DSP_R_X9Y20_DSP48_X0Y8_P1;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_O = LIOB33_X0Y13_IOB_X0Y13_I;
  assign RIOI3_X43Y25_ILOGIC_X1Y26_O = RIOB33_X43Y25_IOB_X1Y26_I;
  assign RIOI3_X43Y39_ILOGIC_X1Y40_O = RIOB33_X43Y39_IOB_X1Y40_I;
  assign RIOI3_X43Y39_ILOGIC_X1Y39_O = RIOB33_X43Y39_IOB_X1Y39_I;
  assign RIOI3_X43Y45_ILOGIC_X1Y46_O = RIOB33_X43Y45_IOB_X1Y46_I;
  assign RIOI3_X43Y45_ILOGIC_X1Y45_O = RIOB33_X43Y45_IOB_X1Y45_I;
  assign RIOI3_X43Y47_ILOGIC_X1Y48_O = RIOB33_X43Y47_IOB_X1Y48_I;
  assign RIOI3_X43Y47_ILOGIC_X1Y47_O = RIOB33_X43Y47_IOB_X1Y47_I;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_OQ = DSP_R_X9Y20_DSP48_X0Y8_P14;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_TQ = 1'b1;
  assign RIOI3_X43Y75_OLOGIC_X1Y76_OQ = DSP_R_X9Y20_DSP48_X0Y8_P13;
  assign RIOI3_X43Y75_OLOGIC_X1Y76_TQ = 1'b1;
  assign RIOI3_X43Y75_OLOGIC_X1Y75_OQ = DSP_R_X9Y20_DSP48_X0Y8_P12;
  assign RIOI3_X43Y75_OLOGIC_X1Y75_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_OQ = DSP_R_X9Y20_DSP48_X0Y8_P11;
  assign RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y44_O = RIOB33_X43Y43_IOB_X1Y44_I;
  assign RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y43_O = RIOB33_X43Y43_IOB_X1Y43_I;
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_OQ = DSP_R_X9Y20_DSP48_X0Y8_P9;
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_OQ = DSP_R_X9Y20_DSP48_X0Y8_P10;
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_OQ = DSP_R_X9Y20_DSP48_X0Y8_P15;
  assign RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_TQ = 1'b1;
  assign LIOB33_X0Y19_IOB_X0Y20_O = DSP_R_X9Y20_DSP48_X0Y8_P2;
  assign LIOB33_X0Y19_IOB_X0Y19_O = DSP_R_X9Y20_DSP48_X0Y8_P3;
  assign LIOI3_X0Y17_OLOGIC_X0Y18_T1 = 1'b1;
  assign LIOB33_X0Y1_IOB_X0Y2_O = DSP_R_X9Y20_DSP48_X0Y8_P8;
  assign LIOB33_X0Y1_IOB_X0Y1_O = DSP_R_X9Y20_DSP48_X0Y8_P7;
  assign LIOI3_X0Y9_ILOGIC_X0Y10_D = LIOB33_X0Y9_IOB_X0Y10_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y9_D = LIOB33_X0Y9_IOB_X0Y9_I;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_D1 = DSP_R_X9Y20_DSP48_X0Y8_P14;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_T1 = 1'b1;
  assign RIOI3_X43Y47_ILOGIC_X1Y48_D = RIOB33_X43Y47_IOB_X1Y48_I;
  assign RIOI3_X43Y47_ILOGIC_X1Y47_D = RIOB33_X43Y47_IOB_X1Y47_I;
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_T1 = 1'b1;
  assign RIOB33_X43Y75_IOB_X1Y76_O = DSP_R_X9Y20_DSP48_X0Y8_P13;
  assign RIOB33_X43Y75_IOB_X1Y75_O = DSP_R_X9Y20_DSP48_X0Y8_P12;
  assign DSP_R_X9Y20_DSP48_X0Y8_RSTA = LIOB33_X0Y13_IOB_X0Y13_I;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_I = CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O;
  assign DSP_R_X9Y20_DSP48_X0Y8_RSTALUMODE = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_RSTB = LIOB33_X0Y13_IOB_X0Y13_I;
  assign DSP_R_X9Y20_DSP48_X0Y8_RSTC = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_RSTCTRL = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_RSTD = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_RSTINMODE = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_RSTM = LIOB33_X0Y13_IOB_X0Y13_I;
  assign DSP_R_X9Y20_DSP48_X0Y8_RSTP = LIOB33_X0Y13_IOB_X0Y13_I;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_D1 = DSP_R_X9Y20_DSP48_X0Y8_P8;
  assign RIOB33_X43Y37_IOB_X1Y37_O = DSP_R_X9Y20_DSP48_X0Y8_P10;
  assign RIOB33_X43Y37_IOB_X1Y38_O = DSP_R_X9Y20_DSP48_X0Y8_P9;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_T1 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_D1 = DSP_R_X9Y20_DSP48_X0Y8_P7;
  assign RIOI3_X43Y75_OLOGIC_X1Y76_D1 = DSP_R_X9Y20_DSP48_X0Y8_P13;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_T1 = 1'b1;
  assign RIOI3_X43Y75_OLOGIC_X1Y76_T1 = 1'b1;
  assign LIOB33_SING_X0Y0_IOB_X0Y0_O = DSP_R_X9Y20_DSP48_X0Y8_P6;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_T1 = 1'b1;
  assign RIOB33_X43Y61_IOB_X1Y61_O = DSP_R_X9Y20_DSP48_X0Y8_P14;
  assign RIOI3_X43Y75_OLOGIC_X1Y75_D1 = DSP_R_X9Y20_DSP48_X0Y8_P12;
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_D1 = DSP_R_X9Y20_DSP48_X0Y8_P10;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_D1 = DSP_R_X9Y20_DSP48_X0Y8_P6;
  assign RIOI3_X43Y75_OLOGIC_X1Y75_T1 = 1'b1;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y44_D = RIOB33_X43Y43_IOB_X1Y44_I;
  assign RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y43_D = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOB33_X0Y17_IOB_X0Y18_O = DSP_R_X9Y20_DSP48_X0Y8_P4;
  assign DSP_R_X9Y20_DSP48_X0Y8_A0 = LIOB33_X0Y11_IOB_X0Y11_I;
  assign DSP_R_X9Y20_DSP48_X0Y8_A1 = LIOB33_X0Y11_IOB_X0Y12_I;
  assign DSP_R_X9Y20_DSP48_X0Y8_A2 = LIOB33_X0Y9_IOB_X0Y10_I;
  assign DSP_R_X9Y20_DSP48_X0Y8_A3 = LIOB33_X0Y9_IOB_X0Y9_I;
  assign DSP_R_X9Y20_DSP48_X0Y8_A4 = LIOB33_X0Y7_IOB_X0Y7_I;
  assign DSP_R_X9Y20_DSP48_X0Y8_A5 = LIOB33_X0Y7_IOB_X0Y8_I;
  assign DSP_R_X9Y20_DSP48_X0Y8_A6 = LIOB33_X0Y5_IOB_X0Y5_I;
  assign DSP_R_X9Y20_DSP48_X0Y8_A7 = LIOB33_X0Y5_IOB_X0Y6_I;
  assign DSP_R_X9Y20_DSP48_X0Y8_A8 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_A9 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_A10 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_A11 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_A12 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_A13 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_A14 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_A15 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_A16 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_A17 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_A18 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_A19 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_A20 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_A21 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_A22 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_A23 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_A24 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_A25 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_A26 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_A27 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_A28 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_A29 = 1'b0;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_D = LIOB33_X0Y7_IOB_X0Y8_I;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_D = LIOB33_X0Y7_IOB_X0Y7_I;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_D1 = DSP_R_X9Y20_DSP48_X0Y8_P1;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_CE = 1'b1;
  assign LIOI3_X0Y11_ILOGIC_X0Y12_D = LIOB33_X0Y11_IOB_X0Y12_I;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_D1 = DSP_R_X9Y20_DSP48_X0Y8_P11;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign LIOB33_X0Y3_IOB_X0Y3_O = DSP_R_X9Y20_DSP48_X0Y8_P0;
  assign LIOB33_X0Y3_IOB_X0Y4_O = DSP_R_X9Y20_DSP48_X0Y8_P5;
  assign LIOI3_X0Y5_ILOGIC_X0Y6_D = LIOB33_X0Y5_IOB_X0Y6_I;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_D1 = DSP_R_X9Y20_DSP48_X0Y8_P2;
  assign LIOI3_X0Y5_ILOGIC_X0Y5_D = LIOB33_X0Y5_IOB_X0Y5_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_D = LIOB33_X0Y11_IOB_X0Y11_I;
  assign RIOB33_X43Y87_IOB_X1Y87_O = DSP_R_X9Y20_DSP48_X0Y8_P15;
  assign RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_T1 = 1'b1;
  assign RIOB33_X43Y31_IOB_X1Y32_O = DSP_R_X9Y20_DSP48_X0Y8_P11;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_D1 = DSP_R_X9Y20_DSP48_X0Y8_P3;
  assign DSP_R_X9Y20_DSP48_X0Y8_ALUMODE0 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_ALUMODE1 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_ALUMODE2 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_ALUMODE3 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_B0 = RIOB33_X43Y39_IOB_X1Y40_I;
  assign DSP_R_X9Y20_DSP48_X0Y8_B1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign DSP_R_X9Y20_DSP48_X0Y8_B2 = RIOB33_X43Y47_IOB_X1Y47_I;
  assign DSP_R_X9Y20_DSP48_X0Y8_B3 = RIOB33_X43Y45_IOB_X1Y46_I;
  assign DSP_R_X9Y20_DSP48_X0Y8_B4 = RIOB33_X43Y39_IOB_X1Y39_I;
  assign DSP_R_X9Y20_DSP48_X0Y8_B5 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign DSP_R_X9Y20_DSP48_X0Y8_B6 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign DSP_R_X9Y20_DSP48_X0Y8_B7 = RIOB33_X43Y47_IOB_X1Y48_I;
  assign DSP_R_X9Y20_DSP48_X0Y8_B8 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_B9 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_B10 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_B11 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_B12 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_B13 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_B14 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_B15 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_B16 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_B17 = 1'b0;
  assign LIOB33_X0Y43_IOB_X0Y43_O = DSP_R_X9Y20_DSP48_X0Y8_P1;
  assign RIOI3_X43Y25_ILOGIC_X1Y26_D = RIOB33_X43Y25_IOB_X1Y26_I;
  assign RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_D1 = DSP_R_X9Y20_DSP48_X0Y8_P15;
  assign RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_T1 = 1'b1;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_D1 = DSP_R_X9Y20_DSP48_X0Y8_P5;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_D1 = DSP_R_X9Y20_DSP48_X0Y8_P9;
  assign RIOI3_X43Y45_ILOGIC_X1Y46_D = RIOB33_X43Y45_IOB_X1Y46_I;
  assign RIOI3_X43Y45_ILOGIC_X1Y45_D = RIOB33_X43Y45_IOB_X1Y45_I;
  assign DSP_R_X9Y20_DSP48_X0Y8_C0 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C1 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C2 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C3 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C4 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C5 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C6 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C7 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C8 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C9 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C10 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C11 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C12 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C13 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C14 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C15 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C16 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C17 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C18 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C19 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C20 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C21 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C22 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C23 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C24 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C25 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C26 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C27 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C28 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C29 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C30 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C31 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C32 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C33 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C34 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C35 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C36 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C37 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C38 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C39 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C40 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C41 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C42 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C43 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C44 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C45 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C46 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_C47 = 1'b1;
  assign RIOI3_X43Y39_ILOGIC_X1Y40_D = RIOB33_X43Y39_IOB_X1Y40_I;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_D1 = DSP_R_X9Y20_DSP48_X0Y8_P0;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I0 = RIOB33_X43Y25_IOB_X1Y26_I;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_CARRYINSEL0 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_CARRYINSEL1 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_CARRYINSEL2 = 1'b0;
  assign RIOI3_X43Y39_ILOGIC_X1Y39_D = RIOB33_X43Y39_IOB_X1Y39_I;
  assign DSP_R_X9Y20_DSP48_X0Y8_CEA1 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_CEA2 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_CEAD = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_CEALUMODE = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_CEB1 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_CEB2 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_CEC = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_CECARRYIN = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_CECTRL = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_CED = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_CEINMODE = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_CEM = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_CEP = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign DSP_R_X9Y20_DSP48_X0Y8_D0 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D1 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D2 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D3 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D4 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D5 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D6 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D7 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D8 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D9 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D10 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D11 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D12 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D13 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D14 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D15 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D16 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D17 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D18 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D19 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D20 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D21 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D22 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D23 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_D24 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_INMODE0 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_INMODE1 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_INMODE2 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_INMODE3 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_INMODE4 = 1'b0;
  assign DSP_R_X9Y20_DSP48_X0Y8_OPMODE0 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_OPMODE1 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_OPMODE2 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_OPMODE3 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_OPMODE4 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_OPMODE5 = 1'b1;
  assign DSP_R_X9Y20_DSP48_X0Y8_OPMODE6 = 1'b0;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_D = LIOB33_X0Y13_IOB_X0Y13_I;
  assign LIOI3_X0Y17_OLOGIC_X0Y18_D1 = DSP_R_X9Y20_DSP48_X0Y8_P4;
endmodule
